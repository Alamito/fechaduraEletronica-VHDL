library verilog;
use verilog.vl_types.all;
entity comp_todos_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end comp_todos_vlg_check_tst;
