library verilog;
use verilog.vl_types.all;
entity reg16bits_vlg_vec_tst is
end reg16bits_vlg_vec_tst;
