library verilog;
use verilog.vl_types.all;
entity regUser16bits_vlg_vec_tst is
end regUser16bits_vlg_vec_tst;
