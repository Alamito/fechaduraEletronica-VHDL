library verilog;
use verilog.vl_types.all;
entity regUser4bits_vlg_vec_tst is
end regUser4bits_vlg_vec_tst;
