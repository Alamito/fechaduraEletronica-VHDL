library verilog;
use verilog.vl_types.all;
entity cont2bits_vlg_vec_tst is
end cont2bits_vlg_vec_tst;
