library verilog;
use verilog.vl_types.all;
entity decod4x16_vlg_vec_tst is
end decod4x16_vlg_vec_tst;
