library verilog;
use verilog.vl_types.all;
entity btn_Sincrono_vlg_vec_tst is
end btn_Sincrono_vlg_vec_tst;
