library verilog;
use verilog.vl_types.all;
entity reg4bit_user_vlg_vec_tst is
end reg4bit_user_vlg_vec_tst;
