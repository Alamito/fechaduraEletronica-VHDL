library verilog;
use verilog.vl_types.all;
entity decod2x4_vlg_vec_tst is
end decod2x4_vlg_vec_tst;
