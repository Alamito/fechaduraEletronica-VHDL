library verilog;
use verilog.vl_types.all;
entity cont1bit_vlg_vec_tst is
end cont1bit_vlg_vec_tst;
