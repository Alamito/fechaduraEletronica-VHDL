library verilog;
use verilog.vl_types.all;
entity reg4bits_vlg_vec_tst is
end reg4bits_vlg_vec_tst;
