library verilog;
use verilog.vl_types.all;
entity proj_final_16bits_vlg_vec_tst is
end proj_final_16bits_vlg_vec_tst;
