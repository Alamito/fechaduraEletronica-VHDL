library verilog;
use verilog.vl_types.all;
entity reg_decod_vlg_vec_tst is
end reg_decod_vlg_vec_tst;
