library verilog;
use verilog.vl_types.all;
entity Vhdl2_vlg_vec_tst is
end Vhdl2_vlg_vec_tst;
