library verilog;
use verilog.vl_types.all;
entity Ureg4bit_vlg_vec_tst is
end Ureg4bit_vlg_vec_tst;
