library verilog;
use verilog.vl_types.all;
entity decod5x6_vlg_vec_tst is
end decod5x6_vlg_vec_tst;
