library verilog;
use verilog.vl_types.all;
entity display_todos_vlg_vec_tst is
end display_todos_vlg_vec_tst;
