library verilog;
use verilog.vl_types.all;
entity reg1bit_vlg_vec_tst is
end reg1bit_vlg_vec_tst;
