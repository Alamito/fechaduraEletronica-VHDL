library verilog;
use verilog.vl_types.all;
entity display16bits_todos_vlg_vec_tst is
end display16bits_todos_vlg_vec_tst;
