library verilog;
use verilog.vl_types.all;
entity reg1bit_vlg_check_tst is
    port(
        out_reg         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end reg1bit_vlg_check_tst;
